/// I2C custom soft core demo
/// @author Daniel Casner <www.danielcasner.org>

module i2c_softcore (
  input reset,
  input clk
  );
